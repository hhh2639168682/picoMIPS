
//opcodes

`define ADD  4'b0000

`define ADDI 4'b0001

`define MUL 4'b0010

`define SUB 4'b0011

`define HOLD 4'b0100


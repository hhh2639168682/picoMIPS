//-----------------------------------------------------
// File Name   : alucodes.sv
// Function    : pMIPS ALU funcRon code definiRons 
// Version: 1,  only 2 funcs
// Author:  hh2u22
// Last rev. 10/04/23
//-----------------------------------------------------
`define RADD 4'b0000
`define RMUL 4'b0001
`define RSUB 4'b0010